module bram11 (clk, we, re, waddr, raddr, wdi, rdo);
    // define RAMinitFile "./init.dat"
    parameter ADDR_WIDTH = 12;
    parameter SIZE = 11;
    parameter BIT_WIDTH = 32;
    input                          clk;
    input                          we, re;
    input [ADDR_WIDTH-1:0]         waddr, raddr;
    input [BIT_WIDTH-1:0]          wdi;
    output reg [BIT_WIDTH-1:0]     rdo;
    reg [BIT_WIDTH-1:0] RAM [SIZE-1:0];
    // initial $readmemh(RAMinitFile, RAM);

    always @(posedge clk)begin
        if(re) rdo <= RAM[raddr>>2];
    end

    always @(posedge clk)begin
        if(we) RAM[waddr>>2] <= wdi;
    end

endmodule